/*
 * @Author: WenJiaBao-2022E8020282071
 * @Date: 2022-10-30 15:55:46
 * @LastEditTime: 2022-10-30 15:58:40
 * @Description: 
 * 
 * Copyright (c) 2022 by WenJiaBao wenjiabao0919@163.com, All Rights Reserved. 
 */
module ysyx_22050058_mul(
    input   clk,
    input   rst,
    
);